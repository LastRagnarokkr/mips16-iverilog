module pc_add(	input[12:0] a, b,
						output[12:0] sum
						);
	assign sum = a + b;
endmodule